// bit field of register CMD
localparam CMD_START = (1 << 0);
localparam CMD_WRITE = (1 << 1);
localparam CMD_READ  = (1 << 2);
localparam CMD_TXACK = (1 << 3);
localparam CMD_STOP  = (1 << 4);
